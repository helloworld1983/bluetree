
module wr_pattern(clk, rst_n, EN, ADDR, DATA);
    input   clk;
    input   rst_n;
    input   EN;
    input   [7:0] ADDR;
    output reg [33:0] DATA;

always @(posedge clk) begin
    if (EN)
        case (ADDR)
8'h0: DATA <= 34'h290000100;
8'h1: DATA <= 34'h3c0000014;
8'h2: DATA <= 34'h290000000;
8'h3: DATA <= 34'h300000040;
8'h4: DATA <= 34'h290000004;
8'h5: DATA <= 34'h300104040;
8'h6: DATA <= 34'h290000008;
8'h7: DATA <= 34'h300208040;
8'h8: DATA <= 34'h29000000c;
8'h9: DATA <= 34'h30030c040;
8'ha: DATA <= 34'h180001fff;
8'hb: DATA <= 34'h182000008;
8'hc: DATA <= 34'h1840003f0;
8'hd: DATA <= 34'h186000007;
8'he: DATA <= 34'h18800000f;
8'hf: DATA <= 34'h18a000002;
8'h10: DATA <= 34'h18c000002;
8'h11: DATA <= 34'h18e00000c;
8'h12: DATA <= 34'h190000618;
8'h13: DATA <= 34'h100000000;
8'h14: DATA <= 34'h120000002;
8'h15: DATA <= 34'h280001230;
8'h16: DATA <= 34'h3abcdabcd;
8'h17: DATA <= 34'h280002340;
8'h18: DATA <= 34'h312341234;
8'h19: DATA <= 34'h0;
8'h1a: DATA <= 34'h0;
8'h1b: DATA <= 34'h0;
8'h1c: DATA <= 34'h0;
8'h1d: DATA <= 34'h0;
8'h1e: DATA <= 34'h0;
8'h1f: DATA <= 34'h0;
8'h20: DATA <= 34'h0;
8'h21: DATA <= 34'h0;
8'h22: DATA <= 34'h0;
8'h23: DATA <= 34'h0;
8'h24: DATA <= 34'h0;
8'h25: DATA <= 34'h0;
8'h26: DATA <= 34'h0;
8'h27: DATA <= 34'h0;
8'h28: DATA <= 34'h0;
8'h29: DATA <= 34'h0;
8'h2a: DATA <= 34'h0;
8'h2b: DATA <= 34'h0;
8'h2c: DATA <= 34'h0;
8'h2d: DATA <= 34'h0;
8'h2e: DATA <= 34'h0;
8'h2f: DATA <= 34'h0;
8'h30: DATA <= 34'h0;
8'h31: DATA <= 34'h0;
8'h32: DATA <= 34'h0;
8'h33: DATA <= 34'h0;
8'h34: DATA <= 34'h0;
8'h35: DATA <= 34'h0;
8'h36: DATA <= 34'h0;
8'h37: DATA <= 34'h0;
8'h38: DATA <= 34'h0;
8'h39: DATA <= 34'h0;
8'h3a: DATA <= 34'h0;
8'h3b: DATA <= 34'h0;
8'h3c: DATA <= 34'h0;
8'h3d: DATA <= 34'h0;
8'h3e: DATA <= 34'h0;
8'h3f: DATA <= 34'h0;
8'h40: DATA <= 34'h0;
8'h41: DATA <= 34'h0;
8'h42: DATA <= 34'h0;
8'h43: DATA <= 34'h0;
8'h44: DATA <= 34'h0;
8'h45: DATA <= 34'h0;
8'h46: DATA <= 34'h0;
8'h47: DATA <= 34'h0;
8'h48: DATA <= 34'h0;
8'h49: DATA <= 34'h0;
8'h4a: DATA <= 34'h0;
8'h4b: DATA <= 34'h0;
8'h4c: DATA <= 34'h0;
8'h4d: DATA <= 34'h0;
8'h4e: DATA <= 34'h0;
8'h4f: DATA <= 34'h0;
8'h50: DATA <= 34'h0;
8'h51: DATA <= 34'h0;
8'h52: DATA <= 34'h0;
8'h53: DATA <= 34'h0;
8'h54: DATA <= 34'h0;
8'h55: DATA <= 34'h0;
8'h56: DATA <= 34'h0;
8'h57: DATA <= 34'h0;
8'h58: DATA <= 34'h0;
8'h59: DATA <= 34'h0;
8'h5a: DATA <= 34'h0;
8'h5b: DATA <= 34'h0;
8'h5c: DATA <= 34'h0;
8'h5d: DATA <= 34'h0;
8'h5e: DATA <= 34'h0;
8'h5f: DATA <= 34'h0;
8'h60: DATA <= 34'h0;
8'h61: DATA <= 34'h0;
8'h62: DATA <= 34'h0;
8'h63: DATA <= 34'h0;
8'h64: DATA <= 34'h0;
8'h65: DATA <= 34'h0;
8'h66: DATA <= 34'h0;
8'h67: DATA <= 34'h0;
8'h68: DATA <= 34'h0;
8'h69: DATA <= 34'h0;
8'h6a: DATA <= 34'h0;
8'h6b: DATA <= 34'h0;
8'h6c: DATA <= 34'h0;
8'h6d: DATA <= 34'h0;
8'h6e: DATA <= 34'h0;
8'h6f: DATA <= 34'h0;
8'h70: DATA <= 34'h0;
8'h71: DATA <= 34'h0;
8'h72: DATA <= 34'h0;
8'h73: DATA <= 34'h0;
8'h74: DATA <= 34'h0;
8'h75: DATA <= 34'h0;
8'h76: DATA <= 34'h0;
8'h77: DATA <= 34'h0;
8'h78: DATA <= 34'h0;
8'h79: DATA <= 34'h0;
8'h7a: DATA <= 34'h0;
8'h7b: DATA <= 34'h0;
8'h7c: DATA <= 34'h0;
8'h7d: DATA <= 34'h0;
8'h7e: DATA <= 34'h0;
8'h7f: DATA <= 34'h0;
8'h80: DATA <= 34'h0;
8'h81: DATA <= 34'h0;
8'h82: DATA <= 34'h0;
8'h83: DATA <= 34'h0;
8'h84: DATA <= 34'h0;
8'h85: DATA <= 34'h0;
8'h86: DATA <= 34'h0;
8'h87: DATA <= 34'h0;
8'h88: DATA <= 34'h0;
8'h89: DATA <= 34'h0;
8'h8a: DATA <= 34'h0;
8'h8b: DATA <= 34'h0;
8'h8c: DATA <= 34'h0;
8'h8d: DATA <= 34'h0;
8'h8e: DATA <= 34'h0;
8'h8f: DATA <= 34'h0;
8'h90: DATA <= 34'h0;
8'h91: DATA <= 34'h0;
8'h92: DATA <= 34'h0;
8'h93: DATA <= 34'h0;
8'h94: DATA <= 34'h0;
8'h95: DATA <= 34'h0;
8'h96: DATA <= 34'h0;
8'h97: DATA <= 34'h0;
8'h98: DATA <= 34'h0;
8'h99: DATA <= 34'h0;
8'h9a: DATA <= 34'h0;
8'h9b: DATA <= 34'h0;
8'h9c: DATA <= 34'h0;
8'h9d: DATA <= 34'h0;
8'h9e: DATA <= 34'h0;
8'h9f: DATA <= 34'h0;
8'ha0: DATA <= 34'h0;
8'ha1: DATA <= 34'h0;
8'ha2: DATA <= 34'h0;
8'ha3: DATA <= 34'h0;
8'ha4: DATA <= 34'h0;
8'ha5: DATA <= 34'h0;
8'ha6: DATA <= 34'h0;
8'ha7: DATA <= 34'h0;
8'ha8: DATA <= 34'h0;
8'ha9: DATA <= 34'h0;
8'haa: DATA <= 34'h0;
8'hab: DATA <= 34'h0;
8'hac: DATA <= 34'h0;
8'had: DATA <= 34'h0;
8'hae: DATA <= 34'h0;
8'haf: DATA <= 34'h0;
8'hb0: DATA <= 34'h0;
8'hb1: DATA <= 34'h0;
8'hb2: DATA <= 34'h0;
8'hb3: DATA <= 34'h0;
8'hb4: DATA <= 34'h0;
8'hb5: DATA <= 34'h0;
8'hb6: DATA <= 34'h0;
8'hb7: DATA <= 34'h0;
8'hb8: DATA <= 34'h0;
8'hb9: DATA <= 34'h0;
8'hba: DATA <= 34'h0;
8'hbb: DATA <= 34'h0;
8'hbc: DATA <= 34'h0;
8'hbd: DATA <= 34'h0;
8'hbe: DATA <= 34'h0;
8'hbf: DATA <= 34'h0;
8'hc0: DATA <= 34'h0;
8'hc1: DATA <= 34'h0;
8'hc2: DATA <= 34'h0;
8'hc3: DATA <= 34'h0;
8'hc4: DATA <= 34'h0;
8'hc5: DATA <= 34'h0;
8'hc6: DATA <= 34'h0;
8'hc7: DATA <= 34'h0;
8'hc8: DATA <= 34'h0;
8'hc9: DATA <= 34'h0;
8'hca: DATA <= 34'h0;
8'hcb: DATA <= 34'h0;
8'hcc: DATA <= 34'h0;
8'hcd: DATA <= 34'h0;
8'hce: DATA <= 34'h0;
8'hcf: DATA <= 34'h0;
8'hd0: DATA <= 34'h0;
8'hd1: DATA <= 34'h0;
8'hd2: DATA <= 34'h0;
8'hd3: DATA <= 34'h0;
8'hd4: DATA <= 34'h0;
8'hd5: DATA <= 34'h0;
8'hd6: DATA <= 34'h0;
8'hd7: DATA <= 34'h0;
8'hd8: DATA <= 34'h0;
8'hd9: DATA <= 34'h0;
8'hda: DATA <= 34'h0;
8'hdb: DATA <= 34'h0;
8'hdc: DATA <= 34'h0;
8'hdd: DATA <= 34'h0;
8'hde: DATA <= 34'h0;
8'hdf: DATA <= 34'h0;
8'he0: DATA <= 34'h0;
8'he1: DATA <= 34'h0;
8'he2: DATA <= 34'h0;
8'he3: DATA <= 34'h0;
8'he4: DATA <= 34'h0;
8'he5: DATA <= 34'h0;
8'he6: DATA <= 34'h0;
8'he7: DATA <= 34'h0;
8'he8: DATA <= 34'h0;
8'he9: DATA <= 34'h0;
8'hea: DATA <= 34'h0;
8'heb: DATA <= 34'h0;
8'hec: DATA <= 34'h0;
8'hed: DATA <= 34'h0;
8'hee: DATA <= 34'h0;
8'hef: DATA <= 34'h0;
8'hf0: DATA <= 34'h0;
8'hf1: DATA <= 34'h0;
8'hf2: DATA <= 34'h0;
8'hf3: DATA <= 34'h0;
8'hf4: DATA <= 34'h0;
8'hf5: DATA <= 34'h0;
8'hf6: DATA <= 34'h0;
8'hf7: DATA <= 34'h0;
8'hf8: DATA <= 34'h0;
8'hf9: DATA <= 34'h0;
8'hfa: DATA <= 34'h0;
8'hfb: DATA <= 34'h0;
8'hfc: DATA <= 34'h0;
8'hfd: DATA <= 34'h0;
8'hfe: DATA <= 34'h0;
8'hff: DATA <= 34'h0;

        endcase
end
endmodule
